/* testbench para Adder16 */
/* ordem de portas: s, ovfl, a, b */
/* input [15:0] a; input [15:0] b; */
/* output [15:0] s; output ovfl; */

`include "Adder16.v"

`define assert(signal, value) \
    if (signal !== value) \
    begin \
        $display("ASSERTION FAILED in %m: signal != value"); \
        $finish; \
    end else begin \
        $display("Success! %m: signal = value"); \
    end

module tb_Adder16;
    reg [15:0] a;
    reg [15:0] b;
    wire [15:0] s;
    wire ovfl;

    Adder16 mymodule(s, ovfl, a, b);
    
    initial
    begin
        $dumpfile("tb_Adder16.vcd");
        $dumpvars(0, tb_Adder16);

        a = 16'b0000000000000000; b = 16'b0000000000000000; #1;
         `assert(s, 16'b0000000000000000) `assert(ovfl, 1'b0)
        a = 16'b0000100001010001; b = 16'b1101111110110101; #1;
         `assert(s, 16'b1110100000000110) `assert(ovfl, 1'b0)
        a = 16'b0001000111111110; b = 16'b1001111010000011; #1;
         `assert(s, 16'b1011000010000001) `assert(ovfl, 1'b0)
        a = 16'b0001001000000101; b = 16'b1100000111011001; #1;
         `assert(s, 16'b1101001111011110) `assert(ovfl, 1'b0)
        a = 16'b0001110101100111; b = 16'b1110001110001100; #1;
         `assert(s, 16'b0000000011110011) `assert(ovfl, 1'b1)
        a = 16'b0011000010001011; b = 16'b0010101110000001; #1;
         `assert(s, 16'b0101110000001100) `assert(ovfl, 1'b0)
        a = 16'b0011111000001111; b = 16'b0110011010001111; #1;
         `assert(s, 16'b1010010010011110) `assert(ovfl, 1'b0)
        a = 16'b0100000011000000; b = 16'b0010111110100001; #1;
         `assert(s, 16'b0111000001100001) `assert(ovfl, 1'b0)
        a = 16'b0100010010110101; b = 16'b1011101010000000; #1;
         `assert(s, 16'b1111111100110101) `assert(ovfl, 1'b0)
        a = 16'b0101010010110100; b = 16'b1110101011110001; #1;
         `assert(s, 16'b0011111110100101) `assert(ovfl, 1'b1)
        a = 16'b0101111110001110; b = 16'b1101100000001011; #1;
         `assert(s, 16'b0011011110011001) `assert(ovfl, 1'b1)
        a = 16'b0111100000010101; b = 16'b1001011110000011; #1;
         `assert(s, 16'b0000111110011000) `assert(ovfl, 1'b1)
        a = 16'b0111111001010101; b = 16'b1101101100101110; #1;
         `assert(s, 16'b0101100110000011) `assert(ovfl, 1'b1)
        a = 16'b1000100010001111; b = 16'b1111100100001011; #1;
         `assert(s, 16'b1000000110011010) `assert(ovfl, 1'b1)
        a = 16'b1000100101110111; b = 16'b1101010101001010; #1;
         `assert(s, 16'b0101111011000001) `assert(ovfl, 1'b1)
        a = 16'b1001100101011001; b = 16'b1111010111100001; #1;
         `assert(s, 16'b1000111100111010) `assert(ovfl, 1'b1)
        a = 16'b1010010111111011; b = 16'b1000001000100111; #1;
         `assert(s, 16'b0010100000100010) `assert(ovfl, 1'b1)
        a = 16'b1010100101001100; b = 16'b0001101011001001; #1;
         `assert(s, 16'b1100010000010101) `assert(ovfl, 1'b0)
        a = 16'b1011101110110110; b = 16'b0111000111000011; #1;
         `assert(s, 16'b0010110101111001) `assert(ovfl, 1'b1)
        a = 16'b1011110101011101; b = 16'b1110010110111011; #1;
         `assert(s, 16'b1010001100011000) `assert(ovfl, 1'b1)
        a = 16'b1011110110011000; b = 16'b1000100100010001; #1;
         `assert(s, 16'b0100011010101001) `assert(ovfl, 1'b1)
        a = 16'b1101111011100110; b = 16'b1111100011110100; #1;
         `assert(s, 16'b1101011111011010) `assert(ovfl, 1'b1)
        a = 16'b1110001000100111; b = 16'b1011001000110010; #1;
         `assert(s, 16'b1001010001011001) `assert(ovfl, 1'b1)
        a = 16'b1110110101010011; b = 16'b0101001100001110; #1;
         `assert(s, 16'b0100000001100001) `assert(ovfl, 1'b1)
        a = 16'b1111001010001100; b = 16'b1011110110000011; #1;
         `assert(s, 16'b1011000000001111) `assert(ovfl, 1'b1)
        a = 16'b1111001100100100; b = 16'b1111111101011001; #1;
         `assert(s, 16'b1111001001111101) `assert(ovfl, 1'b1)
        a = 16'b1111010000010001; b = 16'b1101011011110111; #1;
         `assert(s, 16'b1100101100001000) `assert(ovfl, 1'b1)
        a = 16'b1111011101011011; b = 16'b1001001011101010; #1;
         `assert(s, 16'b1000101001000101) `assert(ovfl, 1'b1)
        a = 16'b1111100111001100; b = 16'b1100111001100010; #1;
         `assert(s, 16'b1100100000101110) `assert(ovfl, 1'b1)
        a = 16'b1111111111111111; b = 16'b1111111111111111; #1;
         `assert(s, 16'b1111111111111110) `assert(ovfl, 1'b1)

    end
endmodule